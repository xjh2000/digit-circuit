module lllwbc_p_inverse (
    input [63:0] state,
    output [63:0] state_next);


endmodule // lllwbc_p_inverse