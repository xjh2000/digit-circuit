module lllwbc_p (
    input [63:0] state,
    output [63:0] state_next);


endmodule // lllwbc_p