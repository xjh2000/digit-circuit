module or_gate (input a,
                input b,
                output wire y);
    assign y = a | b;
endmodule //and_gate
