module not_gate (input a,
                input b,
                output wire y);
    assign y = ~a;
endmodule //and_gate
