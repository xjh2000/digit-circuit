module lllwbc_f (
    input [7:0] state,
    output [7:0] state_next);


endmodule // lllwbc_f