module lllwbc_encrypt (
    input clk,
    input [63:0] plain_text,
    input [127:0] key,
    output [63:0] cipher_text);


endmodule // lllwbc_encrypt