module lllwbc_key_schedule (
    input [127:0] key,
    output [63:0] kws[1:0],
    output [31:0] krs[20:0]);


endmodule // lllwbc_key_schedule